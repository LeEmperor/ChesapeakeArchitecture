// Bohdan Purtell
`timescale 1 ns / 1 ps

module testbench_controller_v1();
    logic [5:0] tb_funct7,
    logic [] tb_funct7,
    
